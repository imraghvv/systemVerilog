interface inf(input logic clk, rst);

logic [1:0]a;
logic [1:0]b;
logic [1:0]o;
logic [1:0]bo;
logic [1:0]c;
logic [1:0]result;

endinterface
