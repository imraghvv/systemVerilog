interface inf(input logic clk,reset);
    logic a;
    logic b;
    logic cin;
    logic s; 
    logic cout;
endinterface //FA